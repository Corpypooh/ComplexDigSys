library ieee;
use ieee.std_logic_1164.all;

entity Lab1_3 is
port(
	------------ KEY ------------
	KEY             	:in    	std_logic_vector(1 downto 0);

	------------ SW ------------
	SW              	:in    	std_logic_vector(1 downto 0);

	------------ LED ------------
	LEDR            	:out   	std_logic_vector(9 downto 0)
	);
end Lab1_3;

architecture shift of Lab1_3 is
	component flipflop
	port (
		D, clk, rst, set		: in	std_logic;
		q							: out std_logic);
	end component;
	
	signal clk	 : std_logic;
	signal rst	 : std_logic;
	signal w 	 : std_logic;
	signal z		 : std_logic;
	signal Q_0 	 : std_logic_vector(3 downto 0);
	signal Q_1 	 : std_logic_vector(3 downto 0);
	--Tie hardware inputs to software signals
begin
	clk 	<= KEY(0);
	rst	<= SW(0);
	w		<= SW(1);
	
	--Shift register for 0000 detection
	ZFF0: flipflop PORT MAP (w, clk, rst, '1', Q_0(0));
	ZFF1: flipflop PORT MAP (Q_0(0), clk, rst, '1', Q_0(1));
	ZFF2: flipflop PORT MAP (Q_0(1), clk, rst, '1', Q_0(2));
	ZFF3: flipflop PORT MAP (Q_0(2), clk, rst, '1', Q_0(3));
	
	--Shift register for 1111 detection
	OFF0: flipflop PORT MAP (w, clk, rst, '1', Q_1(0));
	OFF1: flipflop PORT MAP (Q_1(0), clk, rst, '1', Q_1(1));
	OFF2: flipflop PORT MAP (Q_1(1), clk, rst, '1', Q_1(2));
	OFF3: flipflop PORT MAP (Q_1(2), clk, rst, '1', Q_1(3));

	--Outputs to hardware
	z <= ((Q_0(0) NOR '0') AND (Q_0(1) NOR '0') AND (Q_0(2) NOR '0') AND (Q_0(3) NOR '0')) OR 
			((Q_1(0) AND '1') AND (Q_1(1) AND '1') AND (Q_1(2) AND '1') AND (Q_1(3) AND '1'));
	
	LEDR(3 downto 0) <= Q_0(3 downto 0);
	LEDR(7 downto 4) <= NOT Q_1(3 downto 0);
	
	LEDR(9) <= z;
end shift;
